module PWM_control(

    
);

endmodule // PWM_control